/**
 * JTAG Testbench
 * Tests basic JTAG operations including IDCODE read
 */

`timescale 1ns/1ps

module jtag_tb;
    import jtag_dmi_pkg::*;

    // DPI export for C++ integration
    export "DPI-C" function get_verification_status_dpi;

    reg        clk;
    reg        rst_n;

    // 4 Shared Physical I/O Pins
    reg        jtag_pin0_i;      // Pin 0: TCK/TCKC
    reg        jtag_pin1_i;      // Pin 1: TMS/TMSC input
    wire       jtag_pin1_o;      // Pin 1: TMSC output
    wire       jtag_pin1_oen;    // Pin 1: Output enable (active low)
    reg        jtag_pin2_i;      // Pin 2: TDI
    wire       jtag_pin3_o;      // Pin 3: TDO
    wire       jtag_pin3_oen;    // Pin 3: Output enable (active low)
    reg        jtag_trst_n_i;
    reg        mode_select;

    // DMI interface signals
    wire [DMI_ADDR_WIDTH-1:0] dmi_addr;
    wire [DMI_DATA_WIDTH-1:0] dmi_wdata;
    reg  [DMI_DATA_WIDTH-1:0] dmi_rdata;
    dmi_op_e                  dmi_op;
    dmi_resp_e                dmi_resp;
    wire                      dmi_req_valid;
    reg                       dmi_req_ready;

    wire [31:0] idcode;
    wire       active_mode;

    localparam JTAG_IDCODE = 32'h1DEAD3FF;

    // JTAG module path definitions for easier signal access
    `define JTAG_IR_LATCH    dut.ir_reg.ir_latch
    `define JTAG_IR_OUT      dut.ir_reg.ir_out
    `define JTAG_TAP_STATE   dut.tap_ctrl.state

    // Test tracking variables
    integer test_count = 0;
    integer pass_count = 0;
    integer fail_count = 0;

    // Failed test tracking
    parameter MAX_TESTS = 20;
    string failed_tests [MAX_TESTS];
    integer failed_test_numbers [MAX_TESTS];
    integer failed_test_count = 0;

    // Global variable to track verification results from tasks
    logic last_verification_result = 1'b0;

    logic check1 = 1'b0;
    logic check2 = 1'b0;

    // Task to record failed test
    task record_failed_test(input integer test_num, input string test_name);
        if (failed_test_count < MAX_TESTS) begin
            failed_tests[failed_test_count] = test_name;
            failed_test_numbers[failed_test_count] = test_num;
            failed_test_count = failed_test_count + 1;
        end
    endtask

    // Clock generation
    initial begin
        clk = 0;
        forever #5 clk = ~clk;  // 100MHz clock
    end

    // TCK generation (slower clock for JTAG)
    initial begin
        jtag_pin0_i = 0;
        forever #100 jtag_pin0_i = ~jtag_pin0_i;  // 5MHz JTAG clock
    end

    // DUT instantiation
    jtag_top dut (
        .clk              (clk),
        .rst_n            (rst_n),
        .jtag_pin0_i      (jtag_pin0_i),
        .jtag_pin1_i      (jtag_pin1_i),
        .jtag_pin1_o      (jtag_pin1_o),
        .jtag_pin1_oen    (jtag_pin1_oen),
        .jtag_pin2_i      (jtag_pin2_i),
        .jtag_pin3_o      (jtag_pin3_o),
        .jtag_pin3_oen    (jtag_pin3_oen),
        .jtag_trst_n_i    (jtag_trst_n_i),
        .mode_select      (mode_select),
        .dmi_addr         (dmi_addr),
        .dmi_wdata        (dmi_wdata),
        .dmi_rdata        (dmi_rdata),
        .dmi_op           (dmi_op),
        .dmi_resp         (dmi_resp),
        .dmi_req_valid    (dmi_req_valid),
        .dmi_req_ready    (dmi_req_ready),
        .idcode           (idcode),
        .active_mode      (active_mode)
    );

    // DMI response logic - simple auto-response for testing
    // Returns predictable test patterns based on DMI address to verify
    // proper DMI read operations. Each address returns a unique 32-bit pattern
    // to allow validation of address decoding and data path integrity.
    // This matches the pattern implementation in jtag_vpi_top.sv.
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            dmi_rdata <= 0;
            dmi_resp <= DMI_RESP_SUCCESS;
            dmi_req_ready <= 1'b1;
        end else begin
            dmi_req_ready <= 1'b1;  // Always ready
            dmi_resp <= DMI_RESP_SUCCESS;
            if (dmi_req_valid) begin
                // Return predictable test patterns based on address
                case (dmi_addr)
                    7'h00: dmi_rdata <= 32'hA5A5A5A5;            // Pattern 0
                    7'h01: dmi_rdata <= 32'hAA55AA55;            // Pattern 1
                    7'h02: dmi_rdata <= 32'h55AA55AA;            // Pattern 2 - Used by Test 10
                    7'h03: dmi_rdata <= 32'hFF00FF00;            // Pattern 3
                    7'h04: dmi_rdata <= 32'h00FF00FF;            // Pattern 4
                    7'h05: dmi_rdata <= 32'hACACACAC;            // Pattern 5 - Used by Test 10
                    default: dmi_rdata <= {dmi_addr, dmi_addr, dmi_addr, dmi_addr, 4'h0};  // Address-based pattern
                endcase
            end
        end
    end

    // Test sequence
    initial begin
        // Initialization
        rst_n = 0;
        mode_select = 0;      // Standard JTAG mode
        jtag_pin0_i = 0;
        jtag_pin1_i = 0;
        jtag_pin2_i = 0;
        jtag_trst_n_i = 0;    // Assert reset initially
        dmi_rdata = 0;
        dmi_resp = DMI_RESP_SUCCESS;
        dmi_req_ready = 1;

        #200 rst_n = 1;
        #100 jtag_trst_n_i = 1;  // Release JTAG reset

        $display("=== JTAG Testbench Started ===");
        $display("Time: %0t, Active Mode: %s", $time, active_mode ? "cJTAG" : "JTAG");

        // Test 1: Reset TAP controller
        $display("\nTest 1: TAP Controller Reset");
        test_count = test_count + 1;
        reset_tap();
        read_idcode_with_check(32'h1DEAD3FF);
        if (last_verification_result) begin
            $display("  ✓ TAP reset verification PASSED - IDCODE verification successful");
            pass_count = pass_count + 1;
        end else begin
            $display("  ✗ TAP reset verification FAILED - IDCODE verification failed");
            fail_count = fail_count + 1;
            record_failed_test(1, "TAP Controller Reset");
        end
        #500;

        // Test 2: Read IDCODE (DR scan via default instruction)
        $display("\nTest 2: Read IDCODE (DR scan)");
        test_count = test_count + 1;
        read_idcode_with_check(32'h1DEAD3FF);
        if (last_verification_result) begin
            pass_count = pass_count + 1;
            $display("    ✓ Test 2 PASSED - IDCODE verification successful");
        end else begin
            fail_count = fail_count + 1;
            record_failed_test(2, "Read IDCODE (DR scan)");
            $display("    ✗ Test 2 FAILED - IDCODE verification failed");
        end
        #500;

        // Test 3: IR Scan - Load BYPASS instruction
        $display("\nTest 3: IR Scan - Load BYPASS");
        test_count = test_count + 1;
        write_ir_with_verify(5'h1F);  // BYPASS instruction (5-bit: 0x1F)
        if (last_verification_result) begin
            pass_count = pass_count + 1;
            $display("    ✓ Test 3 PASSED - BYPASS IR instruction loaded successfully");
        end else begin
            fail_count = fail_count + 1;
            record_failed_test(3, "IR Scan - Load BYPASS instruction");
            $display("    ✗ Test 3 FAILED - BYPASS IR instruction load failed");
        end
        #500;

        // Test 4: DR Scan with BYPASS
        $display("\nTest 4: DR Scan - BYPASS register test");
        test_count = test_count + 1;
        reset_tap();  // Reset TAP to ensure clean state
        write_ir_with_verify(5'h1F);  // Reload BYPASS after reset (5-bit: 0x1F)
        test_bypass();
        if (last_verification_result) begin
            pass_count = pass_count + 1;
            $display("    ✓ Test 4 PASSED - BYPASS register test successful");
        end else begin
            fail_count = fail_count + 1;
            record_failed_test(4, "DR Scan - BYPASS register test");
            $display("    ✗ Test 4 FAILED - BYPASS register test failed");
        end
        #500;

        // Test 5: IR Scan - Load IDCODE instruction
        $display("\nTest 5: IR Scan - Load IDCODE instruction");
        test_count = test_count + 1;
        write_ir_with_verify(5'h01);  // Explicitly load IDCODE instruction
        if (last_verification_result) begin
            pass_count = pass_count + 1;
            $display("    ✓ Test 5 PASSED - IDCODE IR instruction loaded successfully");
        end else begin
            fail_count = fail_count + 1;
            record_failed_test(5, "IR Scan - Load IDCODE instruction");
            $display("    ✗ Test 5 FAILED - IDCODE IR instruction load failed");
        end
        #500;

        // Test 6: DR Scan - Read IDCODE
        $display("\nTest 6: DR Scan - Read IDCODE register");
        test_count = test_count + 1;
        read_dr_32bit_with_verify(32'h1DEAD3FF);
        if (last_verification_result) begin
            pass_count = pass_count + 1;
            $display("    ✓ Test 6 PASSED - IDCODE DR read successful");
        end else begin
            fail_count = fail_count + 1;
            record_failed_test(6, "DR Scan - Read IDCODE register");
            $display("    ✗ Test 6 FAILED - IDCODE DR read failed");
        end
        #500;

        // Test 7: IR Scan - Load DTMCS instruction
        $display("\nTest 7: IR Scan - Load DTMCS instruction");
        test_count = test_count + 1;
        write_ir_with_verify(5'h10);  // DTMCS instruction
        if (last_verification_result) begin
            pass_count = pass_count + 1;
            $display("    ✓ Test 7 PASSED - DTMCS IR instruction loaded successfully");
        end else begin
            fail_count = fail_count + 1;
            record_failed_test(7, "IR Scan - Load DTMCS instruction");
            $display("    ✗ Test 7 FAILED - DTMCS IR instruction load failed");
        end
        #500;

        // Test 8: DR Scan - Read DTMCS register
        $display("\nTest 8: DR Scan - Read DTMCS register");
        test_count = test_count + 1;
        read_dr_32bit_with_verify(32'h00001071);  // Expected DTMCS value (RISC-V Debug Spec v0.13.2 compliant)
        if (last_verification_result) begin
            pass_count = pass_count + 1;
            $display("    ✓ Test 8 PASSED - DTMCS DR read successful");
        end else begin
            fail_count = fail_count + 1;
            record_failed_test(8, "DR Scan - Read DTMCS register");
            $display("    ✗ Test 8 FAILED - DTMCS DR read failed");
        end
        #500;

        // Test 9: IR Scan - Load DMI instruction
        $display("\nTest 9: IR Scan - Load DMI instruction");
        test_count = test_count + 1;
        write_ir_with_verify(5'h11);  // DMI instruction
        if (last_verification_result) begin
            pass_count = pass_count + 1;
            $display("    ✓ Test 9 PASSED - DMI IR instruction loaded successfully");
        end else begin
            fail_count = fail_count + 1;
            record_failed_test(9, "IR Scan - Load DMI instruction");
            $display("    ✗ Test 9 FAILED - DMI IR instruction load failed");
        end
        #500;

        // Test 10: DR Scan - Read DMI register (41 bits)
        $display("\nTest 10: DR Scan - Read DMI register");
        test_count = test_count + 1;
        read_dm_register_with_check(7'h02, 32'h55AA55AA);
        check1 = last_verification_result;
        read_dm_register_with_check(7'h05, 32'hACACACAC);
        check2 = last_verification_result;
        if (check1 && check2) begin
            pass_count = pass_count + 1;
            $display("    ✓ Test 10 PASSED - DMI register read successful");
        end else begin
            fail_count = fail_count + 1;
            record_failed_test(10, "DR Scan - Read DMI register");
            $display("    ✗ Test 10 FAILED - DMI register read failed");
        end
        #500;

        // Test 11: Switch to cJTAG mode and read IDCODE
        $display("\nTest 11: cJTAG Mode - Read IDCODE");
        test_count = test_count + 1;
        test_cjtag_idcode_read();
        if (last_verification_result) begin
            pass_count = pass_count + 1;
            $display("    ✓ Test 11 PASSED - cJTAG IDCODE verification successful");
        end else begin
            fail_count = fail_count + 1;
            record_failed_test(11, "cJTAG Mode - Read IDCODE");
            $display("    ✗ Test 11 FAILED - cJTAG IDCODE verification failed");
        end
        #500;

        // Return to JTAG mode
        $display("\nTest 12: Return to JTAG mode");
        test_count = test_count + 1;
        mode_select = 0;
        $display("Returned to JTAG mode, Active Mode: %s", active_mode ? "cJTAG" : "JTAG");
        // Verify JTAG still works after mode switch
        reset_tap();
        read_idcode_with_check(32'h1DEAD3FF);
        if (last_verification_result) begin
            pass_count = pass_count + 1;
            $display("    ✓ Test 12 PASSED - JTAG mode restored and verified");
        end else begin
            fail_count = fail_count + 1;
            record_failed_test(12, "Return to JTAG mode");
            $display("    ✗ Test 12 FAILED - JTAG mode verification failed");
        end
        #200;

        // Test 13: OScan1 OAC Detection
        $display("\nTest 13: OScan1 OAC Detection and Protocol Activation");
        test_count = test_count + 1;
        test_oscan1_oac_detection();
        if (last_verification_result) begin
            pass_count = pass_count + 1;
            $display("    ✓ Test 13 PASSED - OScan1 OAC detection successful");
        end else begin
            fail_count = fail_count + 1;
            record_failed_test(13, "OScan1 OAC Detection and Protocol Activation");
            $display("    ✗ Test 13 FAILED - OScan1 OAC detection failed");
        end
        #500;

        // Test 14: OScan1 JScan Commands
        $display("\nTest 14: OScan1 JScan Command Processing");
        test_count = test_count + 1;
        test_oscan1_jscan_commands();
        if (last_verification_result) begin
            pass_count = pass_count + 1;
            $display("    ✓ Test 14 PASSED - JScan command processing successful");
        end else begin
            fail_count = fail_count + 1;
            record_failed_test(14, "OScan1 JScan Command Processing");
            $display("    ✗ Test 14 FAILED - JScan command processing failed");
        end
        #500;

        // Test 15: OScan1 SF0 Protocol Testing
        $display("\nTest 15: OScan1 Scanning Format 0 (SF0)");
        test_count = test_count + 1;
        test_oscan1_sf0_protocol();
        if (last_verification_result) begin
            pass_count = pass_count + 1;
            $display("    ✓ Test 15 PASSED - SF0 protocol test successful");
        end else begin
            fail_count = fail_count + 1;
            record_failed_test(15, "OScan1 Scanning Format 0 (SF0)");
            $display("    ✗ Test 15 FAILED - SF0 protocol test failed");
        end
        #500;

        // Test 16: OScan1 Zero Insertion/Deletion
        $display("\nTest 16: OScan1 Zero Stuffing (Bit Stuffing)");
        test_count = test_count + 1;
        test_oscan1_zero_stuffing();
        if (last_verification_result) begin
            pass_count = pass_count + 1;
            $display("    ✓ Test 16 PASSED - Zero stuffing test successful");
        end else begin
            fail_count = fail_count + 1;
            record_failed_test(16, "OScan1 Zero Stuffing (Bit Stuffing)");
            $display("    ✗ Test 16 FAILED - Zero stuffing test failed");
        end
        #500;

        // Test 17: Protocol Switching Stress Test
        $display("\nTest 17: JTAG ↔ cJTAG Protocol Switching");
        test_count = test_count + 1;
        test_protocol_switching();
        if (last_verification_result) begin
            pass_count = pass_count + 1;
            $display("    ✓ Test 17 PASSED - Protocol switching successful");
        end else begin
            fail_count = fail_count + 1;
            record_failed_test(17, "JTAG ↔ cJTAG Protocol Switching");
            $display("    ✗ Test 17 FAILED - Protocol switching failed");
        end
        #500;

        // Test 18: Boundary Conditions Testing
        $display("\nTest 18: Protocol Boundary Conditions");
        test_count = test_count + 1;
        test_boundary_conditions();
        if (last_verification_result) begin
            pass_count = pass_count + 1;
            $display("    ✓ Test 18 PASSED - Boundary conditions test successful");
        end else begin
            fail_count = fail_count + 1;
            record_failed_test(18, "Protocol Boundary Conditions");
            $display("    ✗ Test 18 FAILED - Boundary conditions test failed");
        end
        #500;

        // Test 19: Full cJTAG Protocol Test
        $display("\nTest 19: Full cJTAG Protocol Implementation");
        test_count = test_count + 1;
        test_full_cjtag_protocol();
        if (last_verification_result) begin
            pass_count = pass_count + 1;
            $display("    ✓ Test 19 PASSED - Full cJTAG protocol successful");
        end else begin
            fail_count = fail_count + 1;
            record_failed_test(19, "Full cJTAG Protocol Implementation");
            $display("    ✗ Test 19 FAILED - Full cJTAG protocol failed");
        end
        #1000;

        $display("\n=== Enhanced JTAG Testbench Completed ===");
        $display("Tests completed: %0d total, %0d passed, %0d failed", test_count, pass_count, fail_count);

        if (fail_count == 0) begin
            $display("✓ ALL TESTS PASSED!");
            $display("  - TAP Reset and IDCODE verification: PASSED");
            $display("  - Instruction Register operations: PASSED");
            $display("  - Data Register operations: PASSED");
            $display("  - cJTAG/OScan1 protocol: PASSED");
            $display("  - Protocol switching: PASSED");
            $display("  - Boundary conditions: PASSED");
        end else begin
            $display("✗ %0d TESTS FAILED - Details below:", fail_count);
            $display("\n=== FAILED TEST SUMMARY ===");
            for (integer i = 0; i < failed_test_count; i++) begin
                $display("  Test %0d: %s", failed_test_numbers[i], failed_tests[i]);
            end
            $display("\n=== RECOMMENDATIONS ===");
            $display("  - Check waveform file: jtag_sim.fst");
            $display("  - Review JTAG signal timing and protocol");
            $display("  - Verify IDCODE matches expected value (0x1DEAD3FF)");
            $display("  - Check TAP controller state transitions");
        end

        $display("\n=== TEST COVERAGE ===");
        $display("  ✓ IEEE 1149.1 JTAG Protocol");
        $display("  ✓ IEEE 1149.7 cJTAG OScan1 Protocol");
        $display("  ✓ RISC-V Debug Module Interface (DMI)");
        $display("  ✓ Protocol Mode Switching");
        $display("  ✓ Boundary Condition Testing");
        $display("\n=== PERFORMANCE METRICS ===");
        $display("  Total simulation time: %0t", $time);
        $display("  Pass rate: %0d%% (%0d/%0d)", (pass_count * 100) / test_count, pass_count, test_count);

        if (fail_count > 0) begin
            $display("\n=== SIMULATION FAILED ===");
            $finish(1);  // Exit with error code
        end else begin
            $finish;
        end
    end

    // Timeout
    initial begin
        #1000000;
        $display("ERROR: Testbench timeout!");
        $finish(1);  // Exit with error code
    end

    // DPI function wrapper for C++ access
    // Returns: 0 = passed, 1 = failed, 2 = timeout
    function int get_verification_status_dpi();
        int status;
        // Check for timeout condition first
        if ($time >= 1000000) begin
            status = 2;  // Timeout
        end else if (fail_count > 0) begin
            status = 1;  // Failed
        end else if (pass_count > 0 && test_count > 0) begin
            status = 0;  // Passed (has tests and all passed)
        end else begin
            status = 1;  // No tests completed or unknown state - treat as failed
        end
        return status;
    endfunction

    // Task to reset TAP controller
    task reset_tap();
        integer i;
        begin
            $display("  Resetting TAP controller (5 TMS=1 clocks)");
            jtag_pin1_i = 1;
            for (i = 0; i < 5; i = i + 1) begin
                wait_tck();
            end
            jtag_pin1_i = 0;
            wait_tck();
            $display("  TAP reset complete");
        end
    endtask

    // Task to read IDCODE with proper verification
    task read_idcode_with_check(input [31:0] expected_value);
        integer i;
        logic [31:0] read_data;
        begin
            $display("  Reading and verifying IDCODE register...");

            // Go to Run-Test/Idle
            jtag_pin1_i = 0;
            wait_tck();

            // Select DR path (TMS=1)
            jtag_pin1_i = 1;
            wait_tck();

            // Go to Capture-DR (TMS=0)
            jtag_pin1_i = 0;
            wait_tck();

            // Shift IDCODE (shift 32 bits) - use same method as legacy function
            read_data = 32'h0;
            for (i = 0; i < 32; i = i + 1) begin
                jtag_pin2_i = 1'b0;
                jtag_pin1_i = (i == 31) ? 1 : 0;  // TMS=1 on last bit to exit
                wait_tck();
                // Small delay to ensure TDO is stable
                #1;
                read_data = {jtag_pin3_o, read_data[31:1]};
            end

            $display("    IDCODE Read: 0x%08h", read_data);
            $display("    Expected:    0x%08h", expected_value);

            // Check if IDCODE matches expected value and set global result
            if (read_data == expected_value) begin
                $display("    ✓ IDCODE verification PASSED");
                last_verification_result = 1'b1;
            end else begin
                $display("    ✗ IDCODE verification FAILED");
                last_verification_result = 1'b0;
            end

            // Exit shift state (same as legacy function)
            jtag_pin1_i = 1;
            wait_tck();

            // Update-DR
            jtag_pin1_i = 0;
            wait_tck();
        end
    endtask

    // Task to perform proper cJTAG IDCODE read
    task test_cjtag_idcode_read();
        integer i, j;
        logic [31:0] cjtag_idcode;
        logic [3:0] jscan_cmd;
        logic tms_bit, tdi_bit, tdo_captured;
        logic cjtag_working;
        begin
            $display("  Testing cJTAG IDCODE read via OScan1 protocol...");

            // Switch to cJTAG mode
            mode_select = 1;
            #200;
            $display("    Switched to cJTAG mode, Active Mode: %s", active_mode ? "cJTAG" : "JTAG");

            // Send OAC (16 consecutive edges)
            $display("    Sending OAC sequence...");
            for (i = 0; i < 16; i = i + 1) begin
                jtag_pin0_i = ~jtag_pin0_i;
                #25;
            end
            #100;

            // Send JSCAN_OSCAN_ON command (4 bits = 0x1)
            jscan_cmd = 4'h1;  // JSCAN_OSCAN_ON
            $display("    Sending JSCAN_OSCAN_ON command...");
            for (i = 0; i < 4; i = i + 1) begin
                jtag_pin1_i = jscan_cmd[i];  // Send LSB first
                jtag_pin0_i = 1; #25;
                jtag_pin0_i = 0; #25;
            end
            #200;

            // Perform TAP reset via SF0
            $display("    Resetting TAP via SF0 protocol...");
            for (i = 0; i < 5; i = i + 1) begin
                // SF0: TMS on rising edge, TDI on falling edge
                tms_bit = 1; tdi_bit = 0;  // TMS=1 for reset
                jtag_pin1_i = tms_bit; jtag_pin0_i = 1; #25;
                jtag_pin1_i = tdi_bit; jtag_pin0_i = 0; #25;
            end

            // Go to Run-Test-Idle
            tms_bit = 0; tdi_bit = 0;
            jtag_pin1_i = tms_bit; jtag_pin0_i = 1; #25;
            jtag_pin1_i = tdi_bit; jtag_pin0_i = 0; #25;

            // Go to DR scan for IDCODE (should be default after reset)
            // But let's explicitly load IDCODE instruction first

            // Go to IR scan to load IDCODE instruction
            tms_bit = 1; tdi_bit = 0;  // Select-DR to Select-IR
            jtag_pin1_i = tms_bit; jtag_pin0_i = 1; #25;
            jtag_pin1_i = tdi_bit; jtag_pin0_i = 0; #25;

            // Enter Capture-IR (TMS=0)
            tms_bit = 0; tdi_bit = 0;
            jtag_pin1_i = tms_bit; jtag_pin0_i = 1; #25;
            jtag_pin1_i = tdi_bit; jtag_pin0_i = 0; #25;

            // Shift IDCODE instruction (0x01) - 5 bits
            for (j = 0; j < 5; j = j + 1) begin
                tms_bit = (j == 4) ? 1 : 0;  // Exit on last bit
                tdi_bit = (j == 0) ? 1 : 0;  // Send 0x01 (bit 0 = 1, others = 0)
                jtag_pin1_i = tms_bit; jtag_pin0_i = 1; #25;
                jtag_pin1_i = tdi_bit; jtag_pin0_i = 0; #25;
            end

            // Update-IR (TMS=1 from Exit1-IR)
            tms_bit = 1; tdi_bit = 0;
            jtag_pin1_i = tms_bit; jtag_pin0_i = 1; #25;
            jtag_pin1_i = tdi_bit; jtag_pin0_i = 0; #25;

            // Return to Run-Test-Idle (TMS=0)
            tms_bit = 0; tdi_bit = 0;
            jtag_pin1_i = tms_bit; jtag_pin0_i = 1; #25;
            jtag_pin1_i = tdi_bit; jtag_pin0_i = 0; #25;

            // Now go to DR scan for IDCODE
            tms_bit = 1; tdi_bit = 0;
            jtag_pin1_i = tms_bit; jtag_pin0_i = 1; #25;
            jtag_pin1_i = tdi_bit; jtag_pin0_i = 0; #25;

            // Enter Capture-DR (TMS=0)
            tms_bit = 0; tdi_bit = 0;
            jtag_pin1_i = tms_bit; jtag_pin0_i = 1; #25;
            jtag_pin1_i = tdi_bit; jtag_pin0_i = 0; #25;

            // Shift 32 bits of IDCODE using proper SF0 protocol
            $display("    Shifting IDCODE via SF0...");
            cjtag_idcode = 32'h0;
            cjtag_working = 1'b0;

            for (i = 0; i < 32; i = i + 1) begin
                tms_bit = (i == 31) ? 1 : 0;  // TMS=1 on last bit to exit
                tdi_bit = 0;  // Shift zeros for IDCODE read

                // SF0 Rising edge: send TMS bit
                jtag_pin1_i = tms_bit;
                jtag_pin0_i = 1;
                #25;

                // Wait for potential TDO response (give more time)
                #25;

                // Sample TDO if available (check both output enable and data)
                if (jtag_pin1_oen == 1'b0) begin  // oen is active low
                    tdo_captured = jtag_pin1_o;
                    cjtag_idcode = {tdo_captured, cjtag_idcode[31:1]};  // Shift right (LSB first)
                    cjtag_working = 1'b1;  // We got some activity
                    if (i < 8 || i > 23) begin  // Show first/last 8 bits for debug
                        $display("      IDCODE bit %02d: TMS=%b, TDO=%b (captured)", i, tms_bit, tdo_captured);
                    end
                end else begin
                    // No output, use zero
                    cjtag_idcode = {1'b0, cjtag_idcode[31:1]};  // Shift right with zero
                    if (i < 4) begin  // Show first few bits for debug
                        $display("      IDCODE bit %02d: TMS=%b, TDO=0 (no output)", i, tms_bit);
                    end
                end

                // SF0 Falling edge: send TDI bit
                jtag_pin1_i = tdi_bit;
                jtag_pin0_i = 0;
                #25;
            end

            // Exit to Update-DR
            tms_bit = 1; tdi_bit = 0;
            jtag_pin1_i = tms_bit; jtag_pin0_i = 1; #25;
            jtag_pin1_i = tdi_bit; jtag_pin0_i = 0; #25;

            // Return to Run-Test-Idle
            tms_bit = 0; tdi_bit = 0;
            jtag_pin1_i = tms_bit; jtag_pin0_i = 1; #25;
            jtag_pin1_i = tdi_bit; jtag_pin0_i = 0; #25;

            // Check results
            $display("    cJTAG IDCODE: 0x%08h", cjtag_idcode);
            $display("    Expected:     0x%08h", JTAG_IDCODE);

            // More lenient verification - check if we got valid cJTAG activity
            if (cjtag_idcode == JTAG_IDCODE) begin
                $display("    ✓ cJTAG IDCODE verification PASSED - Exact match");
                last_verification_result = 1'b1;
            end else if (cjtag_working && cjtag_idcode != JTAG_IDCODE) begin
                $display("    ✗ cJTAG IDCODE verification FAILED - Got valid cJTAG response");
                last_verification_result = 1'b0;
            end else if (active_mode) begin
                $display("    ✗ cJTAG mode active but OScan1 protocol not fully functional - FAILED");
                last_verification_result = 1'b0;
            end else begin
                $display("    ✗ cJTAG IDCODE verification FAILED - No proper readback");
                last_verification_result = 1'b0;
            end
        end
    endtask

    // Task to write instruction register with verification
    task write_ir_with_verify(input [4:0] instruction);
        integer i;
        logic [4:0] captured_ir;
        logic [4:0] ir_value;
        logic [4:0] expected_value;
        logic capture_passed;
        logic load_passed;
        begin
            ir_value = instruction[4:0];
            expected_value = 5'h01;  // IR capture always returns 0x01 per IEEE 1149.1
            $display("  Writing and verifying IR: 0x%02h (capture will be: 0x%02h)", instruction, expected_value);

            // Go to Run-Test/Idle
            jtag_pin1_i = 0;
            wait_tck();

            // Select IR path (TMS=1, TMS=1)
            jtag_pin1_i = 1;
            wait_tck();
            jtag_pin1_i = 1;
            wait_tck();

            // Go to Capture-IR (TMS=0)
            jtag_pin1_i = 0;
            wait_tck();

            // Transition from Capture-IR to Shift-IR (TMS=0)
            jtag_pin1_i = 0;
            wait_tck();

            // Now in Shift-IR state - shift all 5 bits with proper timing
            captured_ir = 5'h0;
            for (i = 0; i < 5; i = i + 1) begin
                jtag_pin2_i = ir_value[i];  // Set TDI for this bit
                jtag_pin1_i = (i == 4) ? 1 : 0;  // TMS=1 on last bit to exit
                captured_ir = {jtag_pin3_o, captured_ir[4:1]};
                wait_tck();
            end
            $display("    Captured IR: 0x%02h", captured_ir);

            // Now in Exit1-IR state, go to Update-IR (TMS=1)
            jtag_pin1_i = 1;
            wait_tck();

            // Return to Run-Test/Idle (TMS=0 from Update-IR)
            jtag_pin1_i = 0;
            wait_tck();

            // Stay in Run-Test/Idle for a few cycles to let instruction take effect
            repeat(5) wait_tck();

            $display("    Wrote IR: 0x%02h, Captured IR: 0x%02h", ir_value, captured_ir);

            // Dual verification: IEEE 1149.1 compliance + actual instruction load
            capture_passed = (captured_ir == expected_value);
            load_passed = (`JTAG_IR_LATCH == ir_value);

            if (capture_passed) begin
                $display("    ✓ IR capture verification PASSED - IEEE 1149.1 pattern (0x%02h)", expected_value);
            end else begin
                $display("    ✗ IR capture verification FAILED - captured: 0x%02h, expected: 0x%02h", captured_ir, expected_value);
            end

            if (load_passed) begin
                $display("    ✓ IR load verification PASSED - instruction loaded (0x%02h)", ir_value);
            end else begin
                $display("    ✗ IR load verification FAILED - ir_latch: 0x%02h, expected: 0x%02h",
                         `JTAG_IR_LATCH, ir_value);
            end

            // Both verifications must pass
            last_verification_result = capture_passed && load_passed;

            // Debug info
            $display("    Debug: ir_out=0x%02h, tap_state=0x%h", `JTAG_IR_OUT, `JTAG_TAP_STATE);
        end
    endtask

    // Task to read 32-bit data register with verification
    task read_dr_32bit_with_verify(input [31:0] expected_value);
        integer i;
        logic [31:0] read_data;
        begin
            $display("  Reading and verifying 32-bit DR (expected: 0x%08h)...", expected_value);

            // Start from Run-Test/Idle
            jtag_pin1_i = 0;
            wait_tck();

            // Go to Select-DR (TMS=1)
            jtag_pin1_i = 1;
            wait_tck();

            // Go to Capture-DR (TMS=0)
            jtag_pin1_i = 0;
            wait_tck();

            // Shift-DR state - shift 32 bits, with TMS=1 on the last bit
            read_data = 32'h0;
            for (i = 0; i < 32; i = i + 1) begin
                jtag_pin2_i = 1'b0;
                jtag_pin1_i = (i == 31) ? 1 : 0;  // TMS=1 on last bit to exit
                wait_tck();
                #1;
                read_data = {jtag_pin3_o, read_data[31:1]};
            end

            // Exit shift state
            jtag_pin1_i = 1;
            wait_tck();

            // Update-DR
            jtag_pin1_i = 0;
            wait_tck();

            $display("    DR read: 0x%08h", read_data);

            // Verify the read data
            if (read_data == expected_value) begin
                $display("    ✓ DR verification PASSED");
                last_verification_result = 1'b1;
            end else begin
                $display("    ✗ DR verification FAILED");
                last_verification_result = 1'b0;
            end
        end
    endtask

    // Task to wait for TCK edge
    task wait_tck();
        begin
            wait (jtag_pin0_i == 1);
            wait (jtag_pin0_i == 0);
        end
    endtask

    // Task to test BYPASS register
    task test_bypass();
        integer i;
        logic [7:0] test_pattern;
        logic tdo_bit, expected_tdo;
        integer pass_count_local;
        begin
            $display("  Testing BYPASS register...");
            test_pattern = 8'b10110011;
            pass_count_local = 0;
            expected_tdo = 1'b0;  // Initial bypass register state after Capture-DR

            // Start from Run-Test/Idle
            jtag_pin1_i = 0;
            wait_tck();

            // Go to Select-DR (TMS=1)
            jtag_pin1_i = 1;
            wait_tck();

            // Go to Capture-DR (TMS=0) - this loads 0 into bypass register
            jtag_pin1_i = 0;
            wait_tck();

            // Transition to Shift-DR (TMS=0)
            jtag_pin1_i = 0;
            wait_tck();

            // Shift test pattern through BYPASS - need 9 shifts to verify all 8 bits
            // (1 to get captured value, 8 to push all input bits through)
            $display("    Shifting pattern: 0b%08b", test_pattern);
            for (i = 0; i < 9; i = i + 1) begin
                // For first 8 shifts, send pattern bits; for 9th shift, send 0
                if (i < 8) begin
                    jtag_pin2_i = test_pattern[i];
                end else begin
                    jtag_pin2_i = 1'b0;  // Dummy bit to push last pattern bit out
                end

                if (i < 8) begin
                    jtag_pin1_i = 0;  // Stay in Shift-DR for first 8 bits
                end else begin
                    jtag_pin1_i = 1;  // Exit on 9th bit
                end

                // Clock edge happens here - TDI shifts in, TDO shifts out
                wait_tck();

                // Sample TDO after the clock edge
                #1;
                tdo_bit = jtag_pin3_o;

                // Compare with expected
                if (tdo_bit == expected_tdo) begin
                    pass_count_local = pass_count_local + 1;
                    if (i < 8) begin
                        $display("      Bit %0d: TDI=%0b, TDO=%0b (expected=%0b) ✓", i, test_pattern[i], tdo_bit, expected_tdo);
                    end else begin
                        $display("      Bit %0d: TDI=0 (dummy), TDO=%0b (expected=%0b) ✓", i, tdo_bit, expected_tdo);
                    end
                end else begin
                    if (i < 8) begin
                        $display("      Bit %0d: TDI=%0b, TDO=%0b (expected=%0b) ✗", i, test_pattern[i], tdo_bit, expected_tdo);
                    end else begin
                        $display("      Bit %0d: TDI=0 (dummy), TDO=%0b (expected=%0b) ✗", i, tdo_bit, expected_tdo);
                    end
                end

                // Update expected TDO for next iteration
                if (i < 8) begin
                    expected_tdo = test_pattern[i];
                end else begin
                    expected_tdo = 1'b0;  // After dummy bit
                end
            end

            // Update-DR (TMS=1 from Exit1-DR)
            jtag_pin1_i = 1;
            wait_tck();

            // Return to Run-Test/Idle (TMS=0 from Update-DR)
            jtag_pin1_i = 0;
            wait_tck();

            // Check for 9 correct comparisons (captured 0 + pattern[0:7])
            if (pass_count_local >= 9) begin
                $display("    ✓ BYPASS test PASSED (%0d/9 bits correct)", pass_count_local);
                last_verification_result = 1'b1;
            end else begin
                $display("    ✗ BYPASS test FAILED (%0d/9 bits correct)", pass_count_local);
                last_verification_result = 1'b0;
            end
        end
    endtask

    // Task to read DMI register (41 bits) with proper DMI operation
    task read_dm_register_with_check(input [6:0] address, input [31:0] expected_value);
        integer i;
        logic [40:0] write_data, read_data;
        logic [6:0] dmi_addr_test;
        logic [31:0] dmi_data_test;
        logic [1:0] dmi_op_test;
        begin
            $display("  Reading 41-bit DMI register with proper DMI operation...");

            // Step 1: Write a DMI read command to address 0x11 (DMSTATUS)
            dmi_addr_test = address;        // DMSTATUS register address
            dmi_data_test = expected_value; // DMI Data
            dmi_op_test   = 2'b10;          // DMI read operation (01 = write, 10 = read)

            // Construct 41-bit DMI command: [addr:7][data:32][op:2]
            write_data = {dmi_addr_test, dmi_data_test, dmi_op_test};

            $display("    Step 1: Writing DMI read command (addr=0x%02h, op=read)", dmi_addr_test);

            // Start from Run-Test/Idle
            jtag_pin1_i = 0;
            wait_tck();

            // Go to Select-DR (TMS=1)
            jtag_pin1_i = 1;
            wait_tck();

            // Go to Capture-DR (TMS=0)
            jtag_pin1_i = 0;
            wait_tck();

            // Shift-DR state - shift in the DMI command (41 bits)
            for (i = 0; i < 41; i = i + 1) begin
                jtag_pin2_i = write_data[i];  // Shift in LSB first
                jtag_pin1_i = (i == 40) ? 1 : 0;  // TMS=1 on last bit to exit
                wait_tck();
            end

            // Update-DR (TMS=1 from Exit1-DR)
            jtag_pin1_i = 1;
            wait_tck();

            // Return to Run-Test/Idle (TMS=0 from Update-DR)
            jtag_pin1_i = 0;
            wait_tck();

            // Small delay to let DMI operation process
            repeat(5) wait_tck();

            $display("    Step 2: Reading DMI response...");

            // Step 2: Read back the DMI response
            // Go to Select-DR (TMS=1)
            jtag_pin1_i = 1;
            wait_tck();

            // Go to Capture-DR (TMS=0)
            jtag_pin1_i = 0;
            wait_tck();

            // Shift-DR state - shift out the response (41 bits)
            read_data = 41'h0;
            for (i = 0; i < 41; i = i + 1) begin
                jtag_pin2_i = 1'b0;  // Shift in zeros
                jtag_pin1_i = (i == 40) ? 1 : 0;  // TMS=1 on last bit to exit
                wait_tck();
                read_data = {jtag_pin3_o, read_data[40:1]};
            end

            // Update-DR (TMS=1 from Exit1-DR)
            jtag_pin1_i = 1;
            wait_tck();

            // Return to Run-Test/Idle (TMS=0 from Update-DR)
            jtag_pin1_i = 0;
            wait_tck();

            // Parse DMI response fields
            dmi_op_test = read_data[1:0];
            dmi_data_test = read_data[33:2];
            dmi_addr_test = read_data[40:34];

            $display("    DMI response: 0x%011h", read_data);
            $display("      Address: 0x%02h", dmi_addr_test);
            $display("      Data:    0x%08h", dmi_data_test);
            $display("      Op:      0x%01h", dmi_op_test);

            // Verify we got a proper DMI response:
            // - Address should match what we requested (0x11)
            // - Op should be 0 (success) or 2 (in progress)
            // - Data should be non-zero (DMSTATUS has defined bits)
            if (dmi_addr_test == address && (dmi_op_test == 2'h0 || dmi_op_test == 2'h2) && dmi_data_test == expected_value) begin
                $display("    ✓ DMI register operation successful - proper DMI transaction");
                last_verification_result = 1'b1;
            end else begin
                $display("    ✗ DMI register operation failed");
                last_verification_result = 1'b0;
            end
        end
    endtask

    // ========================================
    // Enhanced Protocol Testing Tasks
    // ========================================

    // Task to test OScan1 OAC (Attention Character) detection
    task test_oscan1_oac_detection();
        integer i;
        logic prev_oscan_active;
        logic [3:0] test_cmd;
        logic [31:0] cjtag_test_idcode;
        logic tms_bit, tdi_bit;
        begin
            $display("  Testing OAC detection (16 consecutive edges)...");

            // Switch to cJTAG mode first
            mode_select = 1;
            #100;

            // Capture initial state before OAC
            prev_oscan_active = 1'b0;  // Assume inactive initially
            if ($test$plusargs("oscan_debug")) begin
                // Monitor internal OScan1 controller state if available
                // This would require exposing internal signals in testbench
                $display("    Initial OScan1 state: inactive");
            end

            // Generate 16 consecutive edges on TCKC (jtag_pin0_i)
            $display("    Generating OAC sequence...");
            for (i = 0; i < 16; i = i + 1) begin
                jtag_pin0_i = ~jtag_pin0_i;
                #50; // 50ns edge spacing
            end

            $display("    OAC sequence completed");

            // Wait for OAC detection processing
            #200;

            // Verify OAC detection by attempting JScan command
            // If OAC was detected, we should be able to send JScan commands
            $display("    Verifying OAC detection by testing JScan response...");

            // Try to send a NOOP JScan command (0xF) and monitor for any response
            test_cmd = 4'hF;  // JSCAN_NOOP
            for (i = 0; i < 4; i = i + 1) begin
                jtag_pin1_i = test_cmd[i];
                jtag_pin0_i = 1; #25;
                jtag_pin0_i = 0; #25;
            end
            #100;

            // Verify OAC detection by attempting to read IDCODE in cJTAG mode
            // This provides actual data verification rather than just sequence completion
            $display("    Verifying OAC detection by attempting IDCODE read in cJTAG mode...");

            cjtag_test_idcode = 32'h0;

            // Try a simple JTAG operation via cJTAG to verify the protocol is active
            // Reset TAP via SF0 protocol
            for (i = 0; i < 5; i = i + 1) begin
                tms_bit = 1; tdi_bit = 0;
                jtag_pin1_i = tms_bit; jtag_pin0_i = 1; #25;
                jtag_pin1_i = tdi_bit; jtag_pin0_i = 0; #25;
            end

            // Go to DR scan for IDCODE (should be default after reset)
            tms_bit = 0; tdi_bit = 0;
            jtag_pin1_i = tms_bit; jtag_pin0_i = 1; #25;
            jtag_pin1_i = tdi_bit; jtag_pin0_i = 0; #25;

            tms_bit = 1; tdi_bit = 0;
            jtag_pin1_i = tms_bit; jtag_pin0_i = 1; #25;
            jtag_pin1_i = tdi_bit; jtag_pin0_i = 0; #25;

            tms_bit = 0; tdi_bit = 0;
            jtag_pin1_i = tms_bit; jtag_pin0_i = 1; #25;
            jtag_pin1_i = tdi_bit; jtag_pin0_i = 0; #25;

            // Try to shift a few bits and see if we get any response
            cjtag_test_idcode = 32'h0;
            for (i = 0; i < 8; i = i + 1) begin  // Just test first 8 bits
                tms_bit = (i == 7) ? 1 : 0;  // Exit on last bit
                tdi_bit = 0;

                jtag_pin1_i = tms_bit; jtag_pin0_i = 1; #25;
                if (jtag_pin1_oen) begin
                    cjtag_test_idcode[i] = jtag_pin1_o;
                end
                jtag_pin1_i = tdi_bit; jtag_pin0_i = 0; #25;
            end

            // Update-DR and return to idle
            tms_bit = 1; tdi_bit = 0;
            jtag_pin1_i = tms_bit; jtag_pin0_i = 1; #25;
            jtag_pin1_i = tdi_bit; jtag_pin0_i = 0; #25;
            tms_bit = 0; tdi_bit = 0;
            jtag_pin1_i = tms_bit; jtag_pin0_i = 1; #25;
            jtag_pin1_i = tdi_bit; jtag_pin0_i = 0; #25;

            // Verify we got some response indicating cJTAG protocol is active
            if (cjtag_test_idcode == JTAG_IDCODE) begin
                $display("    ✓ OAC detection test PASSED - cJTAG protocol response detected");
                last_verification_result = 1'b1;
            end else begin
                $display("    ✗ OAC detection test FAILED - No cJTAG response detected");
                last_verification_result = 1'b0;
            end
        end
    endtask

    // Task to test OScan1 JScan command processing
    task test_oscan1_jscan_commands();
        integer i;
        logic [3:0] jscan_cmd;
        logic [7:0] verification_pattern;
        logic [7:0] sf0_captured_data;
        logic sf0_activity_detected;
        begin
            $display("  Testing JScan command processing...");

            // Ensure we're in cJTAG mode
            mode_select = 1;
            #100;

            // Send OAC first to enter JScan mode
            test_oscan1_oac_detection();
            #100;

            // Send JSCAN_OSCAN_ON command (4 bits = 0x1)
            jscan_cmd = 4'h1;  // JSCAN_OSCAN_ON
            $display("    Sending JSCAN_OSCAN_ON (0x1)...");

            for (i = 0; i < 4; i = i + 1) begin
                // Send bit on TMSC during falling edge of TCKC
                jtag_pin1_i = jscan_cmd[i];  // LSB first
                jtag_pin0_i = 1;
                #25;
                jtag_pin0_i = 0;
                #25;
            end

            #200;

            // Verify JScan command was processed by attempting SF0 operation with actual data verification
            $display("    Verifying JSCAN_OSCAN_ON by testing SF0 response with IDCODE attempt...");

            sf0_captured_data = 8'h0;
            sf0_activity_detected = 1'b0;

            // Try SF0 operation: attempt to read partial IDCODE
            // Reset TAP first
            for (i = 0; i < 5; i = i + 1) begin
                // SF0: TMS=1 on rising edge, TDI=0 on falling edge
                jtag_pin1_i = 1'b1;  // TMS bit (reset)
                jtag_pin0_i = 1; #25;
                jtag_pin1_i = 1'b0;  // TDI bit
                jtag_pin0_i = 0; #25;
            end

            // Go to DR scan (TMS sequence: 0,1,0 to reach Shift-DR)
            // Run-Test-Idle (TMS=0)
            jtag_pin1_i = 1'b0; jtag_pin0_i = 1; #25;
            jtag_pin1_i = 1'b0; jtag_pin0_i = 0; #25;
            // Select-DR (TMS=1)
            jtag_pin1_i = 1'b1; jtag_pin0_i = 1; #25;
            jtag_pin1_i = 1'b0; jtag_pin0_i = 0; #25;
            // Capture-DR (TMS=0)
            jtag_pin1_i = 1'b0; jtag_pin0_i = 1; #25;
            jtag_pin1_i = 1'b0; jtag_pin0_i = 0; #25;

            // Try to shift 8 bits and capture response
            for (i = 0; i < 8; i = i + 1) begin
                // SF0: TMS on rising edge, TDI on falling edge
                jtag_pin1_i = (i == 7) ? 1'b1 : 1'b0;  // TMS bit (exit on last)
                jtag_pin0_i = 1; #25;

                // Check for TDO response
                if (jtag_pin1_oen) begin
                    sf0_captured_data[i] = jtag_pin1_o;
                    sf0_activity_detected = 1'b1;
                    $display("      SF0 TDO captured: bit %0d = %b", i, jtag_pin1_o);
                end

                jtag_pin1_i = 1'b0;  // TDI bit (always 0 for read)
                jtag_pin0_i = 0; #25;
            end

            // Exit to Update-DR
            jtag_pin1_i = 1'b1; jtag_pin0_i = 1; #25;
            jtag_pin1_i = 1'b0; jtag_pin0_i = 0; #25;
            // Return to Run-Test-Idle
            jtag_pin1_i = 1'b0; jtag_pin0_i = 1; #25;
            jtag_pin1_i = 1'b0; jtag_pin0_i = 0; #25;

            // Send JSCAN_OSCAN_OFF to exit
            jscan_cmd = 4'h0;  // JSCAN_OSCAN_OFF
            $display("    Sending JSCAN_OSCAN_OFF (0x0)...");

            test_oscan1_oac_detection();  // OAC sequence

            for (i = 0; i < 4; i = i + 1) begin
                jtag_pin1_i = jscan_cmd[i];
                jtag_pin0_i = 1;
                #25;
                jtag_pin0_i = 0;
                #25;
            end

            #200;
            $display("    ✓ JScan OSCAN_OFF command sent - JScan test completed");

            // Verify JScan command processing based on actual SF0 response
            if (sf0_activity_detected && sf0_captured_data != 8'h0) begin // FIXME
                $display("    ✓ JScan command processing test PASSED - SF0 data captured: 0x%02h", sf0_captured_data);
                last_verification_result = 1'b1;
            end else if (sf0_activity_detected) begin
                $display("    ⚠ JScan command processing test - SF0 activity detected but no data");
                last_verification_result = 1'b0;
            end else begin
                $display("    ✗ JScan command processing test FAILED - No SF0 activity detected");
                last_verification_result = 1'b0;
            end
        end
    endtask

    // Task to test OScan1 Scanning Format 0 (SF0)
    task test_oscan1_sf0_protocol();
        integer i;
        logic tms_bit, tdi_bit;
        logic [7:0] sf0_tdo_captured;
        logic [7:0] sf0_pattern;
        begin
            $display("  Testing SF0 scanning format...");

            // Switch to cJTAG mode and activate OScan1
            mode_select = 1;
            #100;

            // Enter OScan1 mode via OAC + JSCAN_ON
            test_oscan1_oac_detection();
            #100;

            // Send JSCAN_OSCAN_ON
            for (i = 0; i < 4; i = i + 1) begin
                jtag_pin1_i = (i == 0) ? 1 : 0;  // 0x1 = JSCAN_OSCAN_ON, LSB first
                jtag_pin0_i = 1; #25; jtag_pin0_i = 0; #25;
            end
            #100;

            $display("    Testing SF0 bit transfer with TDO capture...");

            // Test SF0 protocol with multiple bits and TDO monitoring
            sf0_pattern = 8'b11010010;  // Test pattern
            sf0_tdo_captured = 8'h0;

            for (i = 0; i < 8; i = i + 1) begin
                tms_bit = sf0_pattern[i];
                tdi_bit = 1'(i % 2);  // Alternating TDI pattern

                // SF0 Rising edge: TMS bit
                jtag_pin1_i = tms_bit;
                jtag_pin0_i = 1;
                #25;

                // Check for TDO response during rising edge
                if (jtag_pin1_oen) begin
                    sf0_tdo_captured[i] = jtag_pin1_o;
                    $display("      SF0 bit %0d: TMS=%b, TDO_captured=%b", i, tms_bit, jtag_pin1_o);
                end else begin
                    $display("      SF0 bit %0d: TMS=%b, TDO_not_active", i, tms_bit);
                end

                // SF0 Falling edge: TDI bit
                jtag_pin1_i = tdi_bit;
                jtag_pin0_i = 0;
                #25;
            end

            $display("    SF0 pattern sent: 0x%02h", sf0_pattern);
            $display("    TDO captured:    0x%02h", sf0_tdo_captured);

            // Verify we captured some response
            if (sf0_tdo_captured == sf0_pattern) begin
                $display("    ✓ SF0 protocol test PASSED - TDO activity matches expected patterns");
                last_verification_result = 1'b1;
            end else begin
                $display("    ✗ SF0 protocol test FAILED - No TDO activity detected");
                last_verification_result = 1'b0;
            end
        end
    endtask

    // Task to test OScan1 zero insertion/deletion (bit stuffing)
    task test_oscan1_zero_stuffing();
        integer i;
        logic [7:0] test_pattern;
        logic [15:0] expected_stuffed;  // Pattern with zero insertions
        logic [15:0] observed_pattern;
        begin
            $display("  Testing zero stuffing (bit stuffing)...");

            mode_select = 1;
            #100;

            // Pattern with 5 consecutive ones (should trigger zero insertion)
            test_pattern = 8'b11111010;  // 5 ones followed by other bits
            expected_stuffed = 16'b1111101000010;  // Expected with zero insertion after 5 ones

            $display("    Sending pattern with 5 consecutive ones: 0x%02h", test_pattern);

            // Send OAC and activate OScan1
            test_oscan1_oac_detection();

            // Send JSCAN_OSCAN_ON
            for (i = 0; i < 4; i = i + 1) begin
                jtag_pin1_i = (i == 0) ? 1 : 0;
                jtag_pin0_i = 1; #25; jtag_pin0_i = 0; #25;
            end
            #100;

            // Send test pattern bit by bit and monitor output
            observed_pattern = 16'h0;
            for (i = 0; i < 8; i = i + 1) begin
                jtag_pin1_i = test_pattern[i];
                jtag_pin0_i = 1; #25;

                // Check if zero stuffing is active (would affect timing)
                if (jtag_pin1_oen) begin
                    observed_pattern[i] = jtag_pin1_o;
                    $display("      Bit %0d: Input=%b, Output=%b", i, test_pattern[i], jtag_pin1_o);
                end

                jtag_pin0_i = 0; #25;
            end

            $display("    Input pattern:     0x%02h", test_pattern);
            $display("    Observed pattern:  0x%04h", observed_pattern);

            // Verify bit stuffing behavior (check for any output activity indicating processing)
            if (observed_pattern != 16'h0 || jtag_pin1_oen) begin
                $display("    ✓ Zero stuffing test PASSED - Pattern processing detected");
                last_verification_result = 1'b1;
            end else begin
                $display("    ✗ Zero stuffing test FAILED - No pattern processing detected");
                last_verification_result = 1'b0;
            end
        end
    endtask

    // Task to test protocol switching between JTAG and cJTAG
    task test_protocol_switching();
        logic [31:0] jtag_idcode_1, jtag_idcode_2, cjtag_response;
        logic jtag_mode_verified, cjtag_mode_verified;
        integer j;
        begin
            $display("  Testing protocol switching JTAG ↔ cJTAG...");

            // Start in JTAG mode
            mode_select = 0;
            #200;
            reset_tap();

            // Verify JTAG mode works (without hardcoded expected value)

            $display("    Verifying initial JTAG mode operation...");
            // Read IDCODE in JTAG mode
            jtag_pin1_i = 1; wait_tck();  // Select DR
            jtag_pin1_i = 0; wait_tck();  // Capture DR
            jtag_idcode_1 = 32'h0;
            for (j = 0; j < 32; j = j + 1) begin
                jtag_pin2_i = 1'b0;
                wait_tck();
                jtag_idcode_1 = {jtag_pin3_o, jtag_idcode_1[31:1]};
            end
            jtag_pin1_i = 1; wait_tck();  // Exit
            jtag_pin1_i = 0; wait_tck();
            jtag_mode_verified = (jtag_idcode_1 == JTAG_IDCODE);  // Must match exact expected IDCODE
            $display("      JTAG mode IDCODE: 0x%08h", jtag_idcode_1);

            $display("    Switching to cJTAG mode...");
            mode_select = 1;
            #200;

            // Test basic cJTAG operation
            test_oscan1_oac_detection();
            cjtag_mode_verified = last_verification_result;  // Use result from cJTAG test
            #200;

            $display("    Switching back to JTAG mode...");
            mode_select = 0;
            #200;
            reset_tap();

            // Verify JTAG mode still works after switching
            $display("    Verifying JTAG mode after switching...");
            jtag_pin1_i = 1; wait_tck();  // Select DR
            jtag_pin1_i = 0; wait_tck();  // Capture DR
            jtag_idcode_2 = 32'h0;
            for (j = 0; j < 32; j = j + 1) begin
                jtag_pin2_i = 1'b0;
                wait_tck();
                jtag_idcode_2 = {jtag_pin3_o, jtag_idcode_2[31:1]};
            end
            jtag_pin1_i = 1; wait_tck();  // Exit
            jtag_pin1_i = 0; wait_tck();
            $display("      JTAG mode IDCODE after switching: 0x%08h", jtag_idcode_2);

            $display("    Testing rapid mode switching...");
            repeat(5) begin
                mode_select = ~mode_select;
                #100;
            end

            // Return to JTAG mode
            mode_select = 0;
            #200;

            // Evaluate overall test result - all conditions must pass for a successful test
            $display("    Evaluation results:");
            $display("      - JTAG mode verified: %s", jtag_mode_verified ? "PASS" : "FAIL");
            $display("      - cJTAG mode verified: %s", cjtag_mode_verified ? "PASS" : "FAIL");
            $display("      - IDCODE consistency: %s", (jtag_idcode_1 == jtag_idcode_2) ? "PASS" : "FAIL");
            $display("      - IDCODE exact match: %s", (jtag_idcode_1 == JTAG_IDCODE && jtag_idcode_2 == JTAG_IDCODE) ? "PASS" : "FAIL");

            // Pass only if all critical conditions are met
            if (jtag_mode_verified && cjtag_mode_verified &&
                (jtag_idcode_1 == jtag_idcode_2) && (jtag_idcode_1 == JTAG_IDCODE)) begin
                $display("    ✓ Protocol switching test PASSED - All modes functional, IDCODE exactly correct");
                last_verification_result = 1'b1;
            end else begin
                $display("    ✗ Protocol switching test FAILED - One or more conditions not met");
                if (!jtag_mode_verified) $display("      → JTAG mode verification failed");
                if (!cjtag_mode_verified) $display("      → cJTAG mode verification failed");
                if (jtag_idcode_1 != jtag_idcode_2) $display("      → IDCODE inconsistent before/after mode switch");
                if (jtag_idcode_1 != JTAG_IDCODE) $display("      → First IDCODE incorrect (got 0x%08h, expected 0x1DEAD3FF)", jtag_idcode_1);
                if (jtag_idcode_2 != JTAG_IDCODE) $display("      → Second IDCODE incorrect (got 0x%08h, expected 0x1DEAD3FF)", jtag_idcode_2);
                last_verification_result = 1'b0;
            end
        end
    endtask

    // Task to test boundary conditions
    task test_boundary_conditions();
        integer i;
        logic [31:0] boundary_idcode;
        begin
            $display("  Testing protocol boundary conditions...");

            // Test 1: Very fast mode switching
            $display("    Test 1: Rapid mode switching (10 cycles)");
            for (i = 0; i < 10; i = i + 1) begin
                mode_select = i[0];  // Alternate between 0 and 1
                #10;  // Very fast switching
            end
            mode_select = 0;  // Return to JTAG
            #100;

            // Verify JTAG still works after rapid switching
            $display("    Verifying JTAG functionality after rapid switching...");
            reset_tap();
            read_idcode_with_check(32'h1DEAD3FF);

            // Test 2: Minimum TCKC period in cJTAG mode
            $display("    Test 2: Minimum TCKC period test");
            mode_select = 1;
            #100;
            repeat(20) begin
                jtag_pin0_i = ~jtag_pin0_i;
                #5;  // Very fast clock
            end
            #100;

            // Verify cJTAG mode can handle fast clocking
            // (Check by attempting OAC detection)
            for (i = 0; i < 16; i = i + 1) begin
                jtag_pin0_i = ~jtag_pin0_i;
                #25;  // Normal speed OAC
            end

            // Test 3: Maximum idle time
            $display("    Test 3: Extended idle periods");
            mode_select = 0;
            #1000;  // Long idle period

            // Verify JTAG still works after long idle
            reset_tap();
            read_idcode_with_check(32'h1DEAD3FF);

            // Test 4: Reset during mode switch
            $display("    Test 4: Reset during mode transition");
            mode_select = 1;
            #50;  // Switch mode
            rst_n = 0;  // Reset during transition
            #100;
            rst_n = 1;
            #100;
            mode_select = 0;  // Return to known state
            #200;

            // Verify recovery after reset during transition
            $display("    Verifying recovery after reset during mode transition...");
            reset_tap();

            // Read IDCODE to verify system recovered
            boundary_idcode = 32'h0;
            jtag_pin1_i = 1; wait_tck();  // Select DR
            jtag_pin1_i = 0; wait_tck();  // Capture DR

            for (i = 0; i < 32; i = i + 1) begin
                jtag_pin2_i = 1'b0;
                wait_tck();
                boundary_idcode = {jtag_pin3_o, boundary_idcode[31:1]};
            end

            jtag_pin1_i = 1; wait_tck();  // Exit
            jtag_pin1_i = 0; wait_tck();

            if (boundary_idcode == JTAG_IDCODE) begin
                $display("    ✓ Boundary conditions test PASSED - System recovered properly");
                last_verification_result = 1'b1;
            end else begin
                $display("    ✗ Boundary conditions test FAILED - System did not recover (IDCODE: 0x%08h)", boundary_idcode);
                last_verification_result = 1'b0;
            end
        end
    endtask

    // Task to test full cJTAG protocol implementation
    task test_full_cjtag_protocol();
        integer i, j;
        logic [31:0] cjtag_idcode;
        logic [3:0] jscan_cmd;
        logic tms_bit, tdi_bit, expected_tdo;
        begin
            $display("  Testing complete cJTAG/OScan1 protocol...");

            // Step 1: Switch to cJTAG mode
            mode_select = 1;
            #200;
            $display("    Step 1: Switched to cJTAG mode (mode_select=1)");

            // Step 2: Send OAC (16 consecutive edges to enter JScan mode)
            $display("    Step 2: Sending OAC sequence (16 consecutive TCKC edges)");
            for (i = 0; i < 16; i = i + 1) begin
                jtag_pin0_i = ~jtag_pin0_i;
                #25;  // 25ns per edge, 16 edges = 400ns total
            end
            #100;  // Allow OAC detection to complete

            // Step 3: Send JScan OSCAN_ON command (4 bits: 0x1 = JSCAN_OSCAN_ON)
            $display("    Step 3: Sending JScan OSCAN_ON command (0x1)");
            jscan_cmd = 4'h1;  // JSCAN_OSCAN_ON

            for (i = 0; i < 4; i = i + 1) begin
                // Send JScan command bit by bit (LSB first)
                jtag_pin1_i = jscan_cmd[i];  // TMSC input

                // TCKC rising edge for command bit
                jtag_pin0_i = 1;
                #25;

                // TCKC falling edge
                jtag_pin0_i = 0;
                #25;

                $display("      JScan bit %0d: %b", i, jscan_cmd[i]);
            end
            #200;  // Allow JScan command processing

            // Step 4: Perform SF0 IDCODE read sequence
            // This involves proper 2-phase SF0 protocol:
            // Phase 1: Send TMS=0, TDI=0 to go to Shift-DR and load IDCODE
            $display("    Step 4: SF0 IDCODE read sequence");

            // First, reset TAP via 5 TMS=1 cycles using SF0 protocol
            $display("      Resetting TAP via SF0 (5 cycles TMS=1)");
            for (i = 0; i < 5; i = i + 1) begin
                // SF0: TMS on rising edge, TDI on falling edge
                tms_bit = 1;  // TMS=1 for reset
                tdi_bit = 0;  // TDI=0 (don't care during reset)

                // Rising edge: TMS bit
                jtag_pin1_i = tms_bit;
                jtag_pin0_i = 1;
                #25;

                // Falling edge: TDI bit
                jtag_pin1_i = tdi_bit;
                jtag_pin0_i = 0;
                #25;

                $display("        TAP reset cycle %0d: TMS=%b, TDI=%b", i+1, tms_bit, tdi_bit);
            end

            // Go to Run-Test-Idle (TMS=0)
            tms_bit = 0; tdi_bit = 0;
            jtag_pin1_i = tms_bit; jtag_pin0_i = 1; #25;
            jtag_pin1_i = tdi_bit; jtag_pin0_i = 0; #25;
            $display("      Entered Run-Test-Idle");

            // Enter Select-DR-Scan (TMS=1)
            tms_bit = 1; tdi_bit = 0;
            jtag_pin1_i = tms_bit; jtag_pin0_i = 1; #25;
            jtag_pin1_i = tdi_bit; jtag_pin0_i = 0; #25;

            // Enter Capture-DR (TMS=0)
            tms_bit = 0; tdi_bit = 0;
            jtag_pin1_i = tms_bit; jtag_pin0_i = 1; #25;
            jtag_pin1_i = tdi_bit; jtag_pin0_i = 0; #25;
            $display("      Entered Capture-DR state for IDCODE");

            // Shift 32 bits of IDCODE using SF0 protocol
            $display("      Shifting 32-bit IDCODE via SF0 protocol");
            cjtag_idcode = 32'h0;

            for (i = 0; i < 32; i = i + 1) begin
                // For IDCODE read, we shift zeros and capture TDO
                tms_bit = (i == 31) ? 1 : 0;  // TMS=1 on last bit to exit
                tdi_bit = 0;  // Shift zeros for IDCODE read

                // SF0 Rising edge: TMS bit
                jtag_pin1_i = tms_bit;
                jtag_pin0_i = 1;
                #25;

                // Sample TDO if available (from TMSC output)
                if (jtag_pin1_oen) begin
                    cjtag_idcode[i] = jtag_pin1_o;  // Capture TDO bit
                end

                // SF0 Falling edge: TDI bit
                jtag_pin1_i = tdi_bit;
                jtag_pin0_i = 0;
                #25;

                if (i < 8 || i > 23) begin  // Show first/last 8 bits
                    $display("        IDCODE bit %02d: TMS=%b, TDI=%b, TDO=%b",
                             i, tms_bit, tdi_bit, jtag_pin1_oen ? jtag_pin1_o : 1'bx);
                end
            end

            // Update-DR (TMS=1 from Exit1-DR)
            tms_bit = 1; tdi_bit = 0;
            jtag_pin1_i = tms_bit; jtag_pin0_i = 1; #25;
            jtag_pin1_i = tdi_bit; jtag_pin0_i = 0; #25;

            // Return to Run-Test-Idle
            tms_bit = 0; tdi_bit = 0;
            jtag_pin1_i = tms_bit; jtag_pin0_i = 1; #25;
            jtag_pin1_i = tdi_bit; jtag_pin0_i = 0; #25;

            $display("      cJTAG IDCODE captured: 0x%08h", cjtag_idcode);
            $display("      Expected IDCODE:       0x%08h", JTAG_IDCODE);

            // Step 5: Exit OScan1 mode via JScan OSCAN_OFF
            $display("    Step 5: Sending JScan OSCAN_OFF command");

            // Send OAC again to re-enter JScan mode
            for (i = 0; i < 16; i = i + 1) begin
                jtag_pin0_i = ~jtag_pin0_i;
                #25;
            end
            #100;

            // Send JSCAN_OSCAN_OFF (0x0)
            jscan_cmd = 4'h0;  // JSCAN_OSCAN_OFF
            for (i = 0; i < 4; i = i + 1) begin
                jtag_pin1_i = jscan_cmd[i];
                jtag_pin0_i = 1; #25;
                jtag_pin0_i = 0; #25;
            end
            #200;

            // Step 6: Return to JTAG mode for verification
            $display("    Step 6: Returning to JTAG mode");
            mode_select = 0;
            #200;

            // Verify JTAG mode still works
            reset_tap();
            read_idcode_with_check(32'h1DEAD3FF);

            // Final evaluation
            if (cjtag_idcode == JTAG_IDCODE) begin
                $display("    ✓ Full cJTAG protocol test PASSED");
                $display("      - OAC sequence: Generated successfully");
                $display("      - JScan commands: OSCAN_ON/OSCAN_OFF sent");
                $display("      - SF0 protocol: TMS/TDI phases executed");
                $display("      - IDCODE read: Attempted via 2-wire interface");
                $display("      - Mode switching: JTAG ↔ cJTAG ↔ JTAG");
                last_verification_result = 1'b1;
            end else begin
                $display("    ✗ Full cJTAG protocol test FAILED");
                $display("      - IDCODE mismatch or zero response");
                last_verification_result = 1'b0;
            end

            $display("    Complete IEEE 1149.7 OScan1 protocol validation finished");
        end
    endtask

endmodule
