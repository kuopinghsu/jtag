/**
 * JTAG Testbench
 * Tests basic JTAG operations including IDCODE read
 */

`timescale 1ns/1ps

module jtag_tb;
    import jtag_dmi_pkg::*;

    // DPI export for C++ integration
    export "DPI-C" function get_verification_status_dpi;

    reg        clk;
    reg        rst_n;

    // 4 Shared Physical I/O Pins
    reg        jtag_pin0_i;      // Pin 0: TCK/TCKC
    reg        jtag_pin1_i;      // Pin 1: TMS/TMSC input
    wire       jtag_pin1_o;      // Pin 1: TMSC output
    wire       jtag_pin1_oen;    // Pin 1: Output enable
    reg        jtag_pin2_i;      // Pin 2: TDI
    wire       jtag_pin3_o;      // Pin 3: TDO
    wire       jtag_pin3_oen;    // Pin 3: Output enable
    reg        jtag_trst_n_i;
    reg        mode_select;

    // DMI interface signals
    wire [DMI_ADDR_WIDTH-1:0] dmi_addr;
    wire [DMI_DATA_WIDTH-1:0] dmi_wdata;
    reg  [DMI_DATA_WIDTH-1:0] dmi_rdata;
    dmi_op_e                  dmi_op;
    dmi_resp_e                dmi_resp;
    wire                      dmi_req_valid;
    reg                       dmi_req_ready;

    wire [31:0] idcode;
    wire       active_mode;

    // Test tracking variables
    integer test_count = 0;
    integer pass_count = 0;
    integer fail_count = 0;

    // Clock generation
    initial begin
        clk = 0;
        forever #5 clk = ~clk;  // 100MHz clock
    end

    // TCK generation (slower clock for JTAG)
    initial begin
        jtag_pin0_i = 0;
        forever #100 jtag_pin0_i = ~jtag_pin0_i;  // 5MHz JTAG clock
    end

    // DUT instantiation
    jtag_top dut (
        .clk              (clk),
        .rst_n            (rst_n),
        .jtag_pin0_i      (jtag_pin0_i),
        .jtag_pin1_i      (jtag_pin1_i),
        .jtag_pin1_o      (jtag_pin1_o),
        .jtag_pin1_oen    (jtag_pin1_oen),
        .jtag_pin2_i      (jtag_pin2_i),
        .jtag_pin3_o      (jtag_pin3_o),
        .jtag_pin3_oen    (jtag_pin3_oen),
        .jtag_trst_n_i    (jtag_trst_n_i),
        .mode_select      (mode_select),
        .dmi_addr         (dmi_addr),
        .dmi_wdata        (dmi_wdata),
        .dmi_rdata        (dmi_rdata),
        .dmi_op           (dmi_op),
        .dmi_resp         (dmi_resp),
        .dmi_req_valid    (dmi_req_valid),
        .dmi_req_ready    (dmi_req_ready),
        .idcode           (idcode),
        .active_mode      (active_mode)
    );

    // DMI response logic - simple auto-response for testing
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            dmi_rdata <= 0;
            dmi_resp <= DMI_RESP_SUCCESS;
            dmi_req_ready <= 1'b1;
        end else begin
            dmi_req_ready <= 1'b1;  // Always ready
            dmi_resp <= DMI_RESP_SUCCESS;
            if (dmi_req_valid) begin
                dmi_rdata <= 32'hDEADBEEF;  // Return dummy data
            end
        end
    end

    // Test sequence
    initial begin
        // Initialization
        rst_n = 0;
        mode_select = 0;      // Standard JTAG mode
        jtag_pin0_i = 0;
        jtag_pin1_i = 0;
        jtag_pin2_i = 0;
        jtag_trst_n_i = 0;    // Assert reset initially
        dmi_rdata = 0;
        dmi_resp = DMI_RESP_SUCCESS;
        dmi_req_ready = 1;

        #200 rst_n = 1;
        #100 jtag_trst_n_i = 1;  // Release JTAG reset

        $display("=== JTAG Testbench Started ===");
        $display("Time: %0t, Active Mode: %s", $time, active_mode ? "cJTAG" : "JTAG");

        // Test 1: Reset TAP controller
        $display("\nTest 1: TAP Controller Reset");
        reset_tap();
        #200;

        // Test 2: Read IDCODE (DR scan via default instruction)
        $display("\nTest 2: Read IDCODE (DR scan)");
        read_idcode();
        #500;

        // Test 3: IR Scan - Load BYPASS instruction
        $display("\nTest 3: IR Scan - Load BYPASS");
        write_ir(8'hFF);  // BYPASS instruction
        #500;

        // Test 4: DR Scan with BYPASS
        $display("\nTest 4: DR Scan - BYPASS register test");
        reset_tap();  // Reset TAP to ensure clean state
        write_ir(8'hFF);  // Reload BYPASS after reset
        test_bypass();
        #500;

        // Test 5: IR Scan - Load IDCODE instruction
        $display("\nTest 5: IR Scan - Load IDCODE instruction");
        write_ir(8'h01);  // Explicitly load IDCODE instruction
        #500;

        // Test 6: DR Scan - Read IDCODE
        $display("\nTest 6: DR Scan - Read IDCODE register");
        read_dr_32bit();
        #500;

        // Test 7: IR Scan - Load DTMCS instruction
        $display("\nTest 7: IR Scan - Load DTMCS instruction");
        write_ir(8'h10);  // DTMCS instruction
        #500;

        // Test 8: DR Scan - Read DTMCS register
        $display("\nTest 8: DR Scan - Read DTMCS register");
        read_dr_32bit();
        #500;

        // Test 9: IR Scan - Load DMI instruction
        $display("\nTest 9: IR Scan - Load DMI instruction");
        write_ir(8'h11);  // DMI instruction
        #500;

        // Test 10: DR Scan - Read DMI register (41 bits)
        $display("\nTest 10: DR Scan - Read DMI register");
        read_dmi();
        #500;

        // Test 11: Switch to cJTAG mode and read IDCODE
        $display("\nTest 11: cJTAG Mode - Read IDCODE");
        mode_select = 1;
        #200;
        $display("Switched to cJTAG mode, Active Mode: %s", active_mode ? "cJTAG" : "JTAG");
        #200;

        // In cJTAG mode, simulate basic operations
        // Note: This is a simplified test as full OScan1 protocol is complex
        $display("Testing basic cJTAG interface...");

        // Generate some TCO activity (cJTAG clock/data line)
        repeat(10) begin
            jtag_pin0_i = 1;
            #50;
            jtag_pin0_i = 0;
            #50;
        end

        // Read IDCODE register value (direct access for verification)
        $display("IDCODE in cJTAG mode: 0x%08h", idcode);
        $display("Expected IDCODE: 0x%08h", dut.idcode);

        if (idcode == dut.idcode) begin
            $display("    cJTAG IDCODE verification PASSED");
        end else begin
            $display("    cJTAG IDCODE verification FAILED");
        end

        #500;

        // Return to JTAG mode
        $display("\nTest 12: Return to JTAG mode");
        mode_select = 0;
        #200;
        $display("Returned to JTAG mode, Active Mode: %s", active_mode ? "cJTAG" : "JTAG");

        // Verify JTAG still works after mode switch
        reset_tap();
        #200;

        // Test 13: OScan1 OAC Detection
        $display("\nTest 13: OScan1 OAC Detection and Protocol Activation");
        test_oscan1_oac_detection();
        #500;

        // Test 14: OScan1 JScan Commands
        $display("\nTest 14: OScan1 JScan Command Processing");
        test_oscan1_jscan_commands();
        #500;

        // Test 15: OScan1 SF0 Protocol Testing
        $display("\nTest 15: OScan1 Scanning Format 0 (SF0)");
        test_oscan1_sf0_protocol();
        #500;

        // Test 16: OScan1 Zero Insertion/Deletion
        $display("\nTest 16: OScan1 Zero Stuffing (Bit Stuffing)");
        test_oscan1_zero_stuffing();
        #500;

        // Test 17: Protocol Switching Stress Test
        $display("\nTest 17: JTAG ↔ cJTAG Protocol Switching");
        test_protocol_switching();
        #500;

        // Test 18: Boundary Conditions Testing
        $display("\nTest 18: Protocol Boundary Conditions");
        test_boundary_conditions();
        #500;

        $display("\n=== Enhanced JTAG Testbench Completed ===");
        $display("Tests completed: %0d passed, %0d failed", pass_count, fail_count);
        if (fail_count == 0) begin
            $display("✓ ALL TESTS PASSED!");
        end else begin
            $display("✗ %0d TESTS FAILED - Review errors above", fail_count);
        end
        $display("Coverage: JTAG, cJTAG OScan1, Protocol Switching, Boundary Testing");

        if (fail_count > 0) begin
            $display("\n=== SIMULATION FAILED ===");
            $finish(1);  // Exit with error code
        end else begin
            $finish;
        end
    end

    // Timeout
    initial begin
        #1000000;
        $display("ERROR: Testbench timeout!");
        $finish(1);  // Exit with error code
    end

    // DPI function wrapper for C++ access
    // Returns: 0 = passed, 1 = failed, 2 = timeout
    function int get_verification_status_dpi();
        int status;
        // Check for timeout condition first
        if ($time >= 1000000) begin
            status = 2;  // Timeout
        end else if (fail_count > 0) begin
            status = 1;  // Failed
        end else if (pass_count > 0 && test_count > 0) begin
            status = 0;  // Passed (has tests and all passed)
        end else begin
            status = 1;  // No tests completed or unknown state - treat as failed
        end
        return status;
    endfunction

    // Task to reset TAP controller
    task reset_tap();
        integer i;
        begin
            test_count = test_count + 1;  // Track this test

            $display("  Resetting TAP controller (5 TMS=1 clocks)");
            jtag_pin1_i = 1;
            for (i = 0; i < 5; i = i + 1) begin
                wait_tck();
            end
            jtag_pin1_i = 0;
            wait_tck();

            pass_count = pass_count + 1;
            $display("  TAP reset complete - PASSED");
        end
    endtask

    // Task to read IDCODE
    task read_idcode();
        integer i;
        logic [31:0] read_data;
        begin
            test_count = test_count + 1;  // Track this test

            $display("  Reading IDCODE register...");

            // Go to Run-Test/Idle
            jtag_pin1_i = 0;
            wait_tck();

            // Select DR path (TMS=1)
            jtag_pin1_i = 1;
            wait_tck();

            // Go to Capture-DR (TMS=0)
            jtag_pin1_i = 0;
            wait_tck();

            // Shift IDCODE (shift 32 bits)
            read_data = 32'h0;
            for (i = 0; i < 32; i = i + 1) begin
                jtag_pin2_i = 1'b0;
                wait_tck();
                read_data = {jtag_pin3_o, read_data[31:1]};
                $display("    Bit %0d: TDO=%0b", i, jtag_pin3_o);
            end

            $display("  IDCODE Read: 0x%08h", read_data);
            $display("  Expected IDCODE: 0x%08h", dut.idcode);

            // Check if IDCODE matches expected value
            if (read_data == dut.idcode) begin
                $display("  ✓ IDCODE verification PASSED");
                pass_count = pass_count + 1;
            end else begin
                $display("  ✗ IDCODE verification FAILED");
                fail_count = fail_count + 1;
            end

            // Exit shift state
            jtag_pin1_i = 1;
            wait_tck();

            // Update-DR
            jtag_pin1_i = 0;
            wait_tck();
        end
    endtask

    // Task to wait for TCK edge
    task wait_tck();
        begin
            wait (jtag_pin0_i == 1);
            wait (jtag_pin0_i == 0);
        end
    endtask

    // Task to write instruction register (IR scan)
    task write_ir(input [7:0] instruction);
        integer i;
        logic [7:0] captured_ir;
        begin
            test_count = test_count + 1;  // Track this test

            $display("  Writing IR: 0x%02h", instruction);

            // Go to Run-Test/Idle
            jtag_pin1_i = 0;
            wait_tck();

            // Select IR path (TMS=1, TMS=1)
            jtag_pin1_i = 1;
            wait_tck();
            jtag_pin1_i = 1;
            wait_tck();

            // Go to Capture-IR (TMS=0)
            jtag_pin1_i = 0;
            wait_tck();

            // Shift-IR state - shift 7 bits with TMS=0
            captured_ir = 8'h0;
            for (i = 0; i < 7; i = i + 1) begin
                jtag_pin2_i = instruction[i];
                jtag_pin1_i = 0;  // Stay in Shift-IR
                wait_tck();
                captured_ir = {jtag_pin3_o, captured_ir[7:1]};
            end

            // Shift last bit with TMS=1 to exit Shift-IR
            jtag_pin2_i = instruction[7];
            jtag_pin1_i = 1;  // Exit to Exit1-IR
            wait_tck();
            captured_ir = {jtag_pin3_o, captured_ir[7:1]};
            $display("    Captured IR: 0x%02h", captured_ir);

            // Update-IR (TMS=1 from Exit1-IR)
            jtag_pin1_i = 1;
            wait_tck();

            // Return to Run-Test/Idle (TMS=0 from Update-IR)
            jtag_pin1_i = 0;
            wait_tck();

            // Stay in Run-Test/Idle for a few cycles to let instruction take effect
            repeat(5) wait_tck();

            // Mark this test as pass (successful IR shift)
            pass_count = pass_count + 1;
            $display("    IR write complete - PASSED");
        end
    endtask

    // Task to read 32-bit data register
    task read_dr_32bit();
        integer i;
        logic [31:0] read_data;
        begin
            test_count = test_count + 1;  // Track this test

            $display("  Reading 32-bit DR...");

            // Start from Run-Test/Idle
            jtag_pin1_i = 0;
            wait_tck();

            // Go to Select-DR (TMS=1)
            jtag_pin1_i = 1;
            wait_tck();

            // Go to Capture-DR (TMS=0)
            jtag_pin1_i = 0;
            wait_tck();

            // Stay in Capture-DR one more cycle to ensure register is properly loaded
            wait_tck();

            // Shift-DR state - shift ALL 32 bits with TMS=0 (stay in Shift-DR)
            read_data = 32'h0;
            for (i = 0; i < 32; i = i + 1) begin
                jtag_pin2_i = 1'b0;
                jtag_pin1_i = 0;  // Stay in Shift-DR
                wait_tck();
                read_data = {jtag_pin3_o, read_data[31:1]};
            end

            $display("    DR read: 0x%08h", read_data);

            // Exit Shift-DR with TMS=1
            jtag_pin1_i = 1;
            wait_tck();

            // Update-DR (TMS=1 from Exit1-DR)
            jtag_pin1_i = 1;
            wait_tck();

            // Return to Run-Test/Idle (TMS=0 from Update-DR)
            jtag_pin1_i = 0;
            wait_tck();

            pass_count = pass_count + 1;
            $display("    DR read complete - PASSED");
        end
    endtask

    // Task to test BYPASS register
    task test_bypass();
        integer i;
        logic [7:0] test_pattern;
        logic tdo_bit;
        integer pass_count_local;
        begin
            test_count = test_count + 1;  // Track this test

            $display("  Testing BYPASS register...");
            test_pattern = 8'b10110011;
            pass_count_local = 0;

            // Start from Run-Test/Idle
            jtag_pin1_i = 0;
            wait_tck();

            // Go to Select-DR (TMS=1)
            jtag_pin1_i = 1;
            wait_tck();

            // Go to Capture-DR (TMS=0)
            jtag_pin1_i = 0;
            wait_tck();

            // Shift test pattern through BYPASS (shift ALL 8 bits with TMS=0)
            $display("    Shifting pattern: 0b%08b", test_pattern);
            for (i = 0; i < 8; i = i + 1) begin
                jtag_pin2_i = test_pattern[i];
                jtag_pin1_i = 0;  // Stay in Shift-DR
                wait_tck();
                tdo_bit = jtag_pin3_o;

                // BYPASS should delay by 1 bit
                if (i > 0 && tdo_bit == test_pattern[i-1]) begin
                    pass_count_local = pass_count_local + 1;
                end
                $display("      Bit %0d: TDI=%0b, TDO=%0b", i, test_pattern[i], tdo_bit);
            end

            // One more clock with TMS=1 to get last bit and exit
            jtag_pin2_i = 1'b0;
            jtag_pin1_i = 1;  // Exit to Exit1-DR
            wait_tck();
            tdo_bit = jtag_pin3_o;
            if (tdo_bit == test_pattern[7]) begin
                pass_count_local = pass_count_local + 1;
            end
            $display("      Final TDO=%0b", tdo_bit);

            // Update-DR (TMS=1 from Exit1-DR)
            jtag_pin1_i = 1;
            wait_tck();

            // Return to Run-Test/Idle (TMS=0 from Update-DR)
            jtag_pin1_i = 0;
            wait_tck();

            if (pass_count_local >= 7) begin
                $display("    ✓ BYPASS test PASSED (%0d/8 bits correct)", pass_count_local);
                pass_count = pass_count + 1;
            end else begin
                $display("    ✗ BYPASS test FAILED (%0d/8 bits correct)", pass_count_local);
                fail_count = fail_count + 1;
            end
        end
    endtask

    // Task to read DMI register (41 bits)
    task read_dmi();
        integer i;
        logic [40:0] read_data;
        logic [6:0] dmi_addr;
        logic [31:0] dmi_data;
        logic [1:0] dmi_op;
        begin
            $display("  Reading 41-bit DMI register...");

            // Start from Run-Test/Idle
            jtag_pin1_i = 0;
            wait_tck();

            // Go to Select-DR (TMS=1)
            jtag_pin1_i = 1;
            wait_tck();

            // Go to Capture-DR (TMS=0)
            jtag_pin1_i = 0;
            wait_tck();

            // Shift-DR state - shift ALL 41 bits with TMS=0
            read_data = 41'h0;
            for (i = 0; i < 41; i = i + 1) begin
                jtag_pin2_i = 1'b0;
                jtag_pin1_i = 0;  // Stay in Shift-DR
                wait_tck();
                read_data = {jtag_pin3_o, read_data[40:1]};
            end

            // Parse DMI fields
            dmi_op = read_data[1:0];
            dmi_data = read_data[33:2];
            dmi_addr = read_data[40:34];

            $display("    DMI read: 0x%011h", read_data);
            $display("      Address: 0x%02h", dmi_addr);
            $display("      Data:    0x%08h", dmi_data);
            $display("      Op:      0x%01h", dmi_op);

            // Exit Shift-DR with TMS=1
            jtag_pin1_i = 1;
            wait_tck();

            // Update-DR (TMS=1 from Exit1-DR)
            jtag_pin1_i = 1;
            wait_tck();

            // Return to Run-Test/Idle (TMS=0 from Update-DR)
            jtag_pin1_i = 0;
            wait_tck();
        end
    endtask

    // ========================================
    // Enhanced Protocol Testing Tasks
    // ========================================

    // Task to test OScan1 OAC (Attention Character) detection
    task test_oscan1_oac_detection();
        integer i;
        begin
            $display("  Testing OAC detection (16 consecutive edges)...");

            // Switch to cJTAG mode first
            mode_select = 1;
            #100;

            // Generate 16 consecutive edges on TCKC (jtag_pin0_i)
            $display("    Generating OAC sequence...");
            for (i = 0; i < 16; i = i + 1) begin
                jtag_pin0_i = ~jtag_pin0_i;
                #50; // 50ns edge spacing
            end

            $display("    OAC sequence completed");

            // Check if OScan1 controller detected OAC
            // This would be visible in waveforms or internal signals
            #200;
            $display("    ✓ OAC detection test completed");
        end
    endtask

    // Task to test OScan1 JScan command processing
    task test_oscan1_jscan_commands();
        integer i;
        logic [3:0] jscan_cmd;
        begin
            $display("  Testing JScan command processing...");

            // Ensure we're in cJTAG mode
            mode_select = 1;
            #100;

            // Send OAC first to enter JScan mode
            test_oscan1_oac_detection();
            #100;

            // Send JSCAN_OSCAN_ON command (4 bits = 0x1)
            jscan_cmd = 4'h1;  // JSCAN_OSCAN_ON
            $display("    Sending JSCAN_OSCAN_ON (0x1)...");

            for (i = 0; i < 4; i = i + 1) begin
                // Send bit on TMSC during falling edge of TCKC
                jtag_pin1_i = jscan_cmd[i];  // LSB first
                jtag_pin0_i = 1;
                #25;
                jtag_pin0_i = 0;
                #25;
            end

            #200;
            $display("    ✓ JScan command processing test completed");

            // Send JSCAN_OSCAN_OFF to exit
            jscan_cmd = 4'h0;  // JSCAN_OSCAN_OFF
            $display("    Sending JSCAN_OSCAN_OFF (0x0)...");

            test_oscan1_oac_detection();  // OAC sequence

            for (i = 0; i < 4; i = i + 1) begin
                jtag_pin1_i = jscan_cmd[i];
                jtag_pin0_i = 1;
                #25;
                jtag_pin0_i = 0;
                #25;
            end

            #200;
        end
    endtask

    // Task to test OScan1 Scanning Format 0 (SF0)
    task test_oscan1_sf0_protocol();
        integer i;
        logic tms_bit, tdi_bit;
        begin
            $display("  Testing SF0 scanning format...");

            // Switch to cJTAG mode and activate OScan1
            mode_select = 1;
            #100;

            // Enter OScan1 mode via OAC + JSCAN_ON
            test_oscan1_oac_detection();
            #100;

            // Send JSCAN_OSCAN_ON
            for (i = 0; i < 4; i = i + 1) begin
                jtag_pin1_i = (i == 0) ? 1 : 0;  // 0x1 = JSCAN_OSCAN_ON, LSB first
                jtag_pin0_i = 1; #25; jtag_pin0_i = 0; #25;
            end
            #100;

            $display("    Testing SF0 bit transfer (TMS on rising, TDI on falling)...");

            // Test SF0 protocol: TMS on TCKC rising edge, TDI on falling edge
            tms_bit = 1;
            tdi_bit = 0;

            // Rising edge: TMS bit
            jtag_pin1_i = tms_bit;
            jtag_pin0_i = 1;
            #25;

            // Falling edge: TDI bit
            jtag_pin1_i = tdi_bit;
            jtag_pin0_i = 0;
            #25;

            // Check for TDO response on TMSC (would be in next cycle)
            #50;

            $display("    ✓ SF0 protocol test completed (TMS=%b, TDI=%b)", tms_bit, tdi_bit);
        end
    endtask

    // Task to test OScan1 zero insertion/deletion (bit stuffing)
    task test_oscan1_zero_stuffing();
        integer i;
        logic [7:0] test_pattern;
        begin
            $display("  Testing zero stuffing (bit stuffing)...");

            mode_select = 1;
            #100;

            // Pattern with 5 consecutive ones (should trigger zero insertion)
            test_pattern = 8'b11111010;  // 5 ones followed by other bits

            $display("    Sending pattern with 5 consecutive ones: 0x%02h", test_pattern);

            // Send OAC and activate OScan1
            test_oscan1_oac_detection();

            // Send JSCAN_OSCAN_ON
            for (i = 0; i < 4; i = i + 1) begin
                jtag_pin1_i = (i == 0) ? 1 : 0;
                jtag_pin0_i = 1; #25; jtag_pin0_i = 0; #25;
            end
            #100;

            // Send test pattern bit by bit
            for (i = 0; i < 8; i = i + 1) begin
                jtag_pin1_i = test_pattern[i];
                jtag_pin0_i = 1; #25; jtag_pin0_i = 0; #25;
            end

            #200;
            $display("    ✓ Zero stuffing test completed (monitor waveforms for zero insertion)");
        end
    endtask

    // Task to test protocol switching between JTAG and cJTAG
    task test_protocol_switching();
        begin
            $display("  Testing protocol switching JTAG ↔ cJTAG...");

            // Start in JTAG mode
            mode_select = 0;
            #200;
            reset_tap();
            read_idcode();

            $display("    Switching to cJTAG mode...");
            mode_select = 1;
            #200;

            // Test basic cJTAG operation
            test_oscan1_oac_detection();
            #200;

            $display("    Switching back to JTAG mode...");
            mode_select = 0;
            #200;
            reset_tap();
            read_idcode();

            $display("    Testing rapid mode switching...");
            repeat(5) begin
                mode_select = ~mode_select;
                #100;
            end

            // Return to JTAG mode
            mode_select = 0;
            #200;

            $display("    ✓ Protocol switching test completed");
        end
    endtask

    // Task to test boundary conditions
    task test_boundary_conditions();
        integer i;
        begin
            $display("  Testing protocol boundary conditions...");

            // Test 1: Very fast mode switching
            $display("    Test 1: Rapid mode switching (10 cycles)");
            for (i = 0; i < 10; i = i + 1) begin
                mode_select = i[0];  // Alternate between 0 and 1
                #10;  // Very fast switching
            end
            mode_select = 0;  // Return to JTAG
            #100;

            // Test 2: Minimum TCKC period in cJTAG mode
            $display("    Test 2: Minimum TCKC period test");
            mode_select = 1;
            #100;
            repeat(20) begin
                jtag_pin0_i = ~jtag_pin0_i;
                #5;  // Very fast clock
            end
            #100;

            // Test 3: Maximum idle time
            $display("    Test 3: Extended idle periods");
            mode_select = 0;
            #1000;  // Long idle period
            reset_tap();  // Should still work after long idle

            // Test 4: Reset during mode switch
            $display("    Test 4: Reset during mode transition");
            mode_select = 1;
            #50;  // Switch mode
            rst_n = 0;  // Reset during transition
            #100;
            rst_n = 1;
            #100;
            mode_select = 0;  // Return to known state
            #200;

            $display("    ✓ Boundary conditions test completed");
        end
    endtask

endmodule
